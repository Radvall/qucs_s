.SUBCKT XFMR 1 2 3 4 RATIO=1
E 5 4 1 2 {RATIO}
F 1 2 VM {RATIO}
VM 5 6
RP 1 2 1MEG
RS 6 3 1U
.ENDS
